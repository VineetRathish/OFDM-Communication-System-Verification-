package ofdm_pkg;

import uvm_pkg::*;
`include "seq_item.sv"
`include "sequence.sv"
`include "sequencer.sv"

`include "encoder.sv"
`include "IFFT.sv"
`include "Slicing.sv"
`include "FFT.sv"
`include "driver.sv"
`include "monitor_dut.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "test.sv"

endpackage 
